module rom(
input clock,
input [11:0]address,
output reg [31:0]q
);

always @ (posedge clock)begin
	/*case(address)
	12'h000    :   q<=32'b00000000000000001110001100110111;
	12'h001    :   q<=32'b00000000100000110000001100010011;
	12'h002    :   q<=32'b00000000000000000001001110110111;
	12'h003    :   q<=32'b00000000011100110010000000100011;
	12'h004    :   q<=32'b00000000000000000000001110110111;
	12'h005    :   q<=32'b11111111000000111000001110010011;
	12'h006    :   q<=32'b00110000010100111001000001110011;
	12'h007    :   q<=32'b00110000000001000110000001110011; 
	12'h008	   :   q<=32'b00001000000000000000001100010011;
	12'h009	   :   q<=32'b00110000010000110010000001110011;
	12'h00a    :   q<=32'b00000000000000000000000000010011;
        12'h00b    :   q<=32'b11111110000000000000111101100011;
	default   :   q<=32'b0; 
endcase
*/

	case(address)
	12'h000	:	q<=32'b11111111110000000000001100010011;
	12'h001 :	q<=32'b00000000000000000000001110010011;
	12'h002	:	q<=32'b00000000011100110000000110100011;
	12'h003 :	q<=32'b00000001110000000000010000010011;
	12'h004 :	q<=32'b00000000100000110000000010100011;
	12'h005 : 	q<=32'b00000000000100000000001110010011;
	12'h006 : 	q<=32'b00000000011100110000000000100011;
	12'h007 :	q<=32'b00000001100000000000010000010011;
	12'h008 : 	q<=32'b00000000100000110000000010100011;
	12'h009 : 	q<=32'b00000001110100000000010000010011;
	12'h00a :	q<=32'b00000000100000110000000010100011;
	12'h00b :	q<=32'b00000110000100000000001110010011;
	12'h00c : 	q<=32'b00000000011100110000000000100011;
	12'h00d : 	q<=32'b00000001100100000000010000010011;
	12'h00e :	q<=32'b00000000100000110000000010100011;
	12'h00f :	q<=32'b00000001110100000000010000010011;
	12'h010:	q<=32'b00000000100000110000000010100011;
	default:	q<=32'b0;
endcase

end

endmodule
